 sequence access_state();
    ( !pselx && !penable) ;
  endsequence:access_state
  