

 package master_package;
import uvm_pkg::*;

`include "apb_master_seq_item.sv"
`include "apb_master_sequencer.sv"
`include "apb_master_base_sequence.sv"
`include "apb_master_driver.sv"
`include "apb_master_monitor.sv"
`include "apb_master_config_agent.sv"
`include "apb_master_agent.sv"
`include "apb_scoreboard.sv"
`include "apb_functional_coverage.sv"
`include "apb_master_environment.sv"
`include "apb_base_test.sv"
`include "apb_test_cases.sv"

endpackage:master_package